//Control module for Multi-cycle CPU
//Sequentially controlled, using State machine and ROM

//File includes
`include "opcodes.v"    //"opcodes.v" includes opcode information for all 23 instructions & ALUOp information
`include "states.v"     //"states.v" includes state encoding information for all 26 states

//GENERAL COMMENTS on variable names
//"r_" prefix indicates that the variable is a reg type
//names in "AaaBbb" format are control signals generated by the control module
//names in "aaa_bbb" format are data bits (num_inst is for debugging purpose)

//Module declaration
module Control(clk, reset_n, opcode, function_code, Halt, PCSource, PCWrite, PCWriteCond, IorD, MemRead, MemWrite, IRWrite, RegDst, MemtoReg, RegWrite, ALUSrcA, ALUSrcB, ALUOp, OutWrite, num_inst);
    input clk;
    input reset_n;
    input [3:0] opcode;
    input [5:0] function_code;

    output Halt;
    output [1:0] PCSource;
    output PCWrite;
    output PCWriteCond;
    output IorD;
    output MemRead;
    output MemWrite;
    output IRWrite;
    output [1:0] RegDst;
    output MemtoReg;
    output RegWrite;
    output ALUSrcA;
    output [1:0] ALUSrcB;
    output [3:0] ALUOp;
    output OutWrite;
    output [15:0] num_inst;

    //Internal reg declaration
    reg [4:0] present_state;
    reg [4:0] next_state;

    //to assign control signals inside always block
    reg r_Halt;
    reg [1:0] r_PCSource;
    reg r_PCWrite;
    reg r_PCWriteCond;
    reg r_IorD;
    reg r_MemRead;
    reg r_MemWrite;
    reg r_IRWrite;
    reg [1:0] r_RegDst;
    reg r_MemtoReg;
    reg r_RegWrite;
    reg r_ALUSrcA;
    reg [1:0] r_ALUSrcB;
    reg [3:0] r_ALUOp;
    reg r_OutWrite;
    reg [`WORD_SIZE-1:0] r_num_inst;
    reg [`WORD_SIZE-1:0] r_next_num_inst;
    
    assign Halt = r_Halt;
    assign PCSource = r_PCSource;
    assign PCWrite = r_PCWrite;
    assign PCWriteCond = r_PCWriteCond;
    assign IorD = r_IorD;
    assign MemRead = r_MemRead;
    assign MemWrite = r_MemWrite;
    assign IRWrite = r_IRWrite;
    assign RegDst = r_RegDst;
    assign MemtoReg = r_MemtoReg;
    assign RegWrite = r_RegWrite;
    assign ALUSrcA = r_ALUSrcA;
    assign ALUSrcB = r_ALUSrcB;
    assign ALUOp = r_ALUOp;
    assign OutWrite = r_OutWrite;

    assign num_inst = r_num_inst;

    //Initial state: IDLE
    initial begin
        present_state <= `IDLE;
        r_num_inst <= 1;
        r_next_num_inst <= 1;
    end

    //State machine:
    //  next state logic &
    //  control signal output (as read from ROM)
    always @(present_state, opcode, function_code) begin
        case(present_state)
            //IDLE Stage (after reset, or initial stage)
            `IDLE: begin next_state <= `IF;
                    r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                    end
            //HALT Stage (after machine halts; staying stage after HLT is met)
            `HALT: begin next_state <= `HALT;
                    r_Halt<=1; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                    end

            //IF Stage
            `IF: begin next_state <= `ID;
                    r_IorD<=0; r_MemRead<=1; r_IRWrite<=1;
                    r_ALUSrcA<=0; r_ALUSrcB<=2; r_ALUOp<=`ALUCODE_ADD;
                    r_PCSource<=0; r_PCWrite<=1; r_PCWriteCond<=0;
                    r_Halt<=0; r_MemWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                    end

            //ID Stage
            `ID: case(opcode)
                    //R-type, I-type arithmetic
                    `OPCODE_R: case(function_code)
                            `FUNC_ADD: begin next_state <= `ADD_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_SUB: begin next_state <= `SUB_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_AND: begin next_state <= `AND_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_ORR: begin next_state <= `ORR_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_NOT: begin next_state <= `NOT_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_TCP: begin next_state <= `TCP_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_SHL: begin next_state <= `SHL_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            `FUNC_SHR: begin next_state <= `SHR_EX;
                                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                        end
                            //JPR
                            `FUNC_JPR: begin next_state <= `IF;
                                    r_PCSource<=2; r_PCWrite<=1; r_PCWriteCond<=0;
                                    r_Halt<=0; r_MemRead<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                                    r_next_num_inst <= r_num_inst + 1;
                                    end
                            //JRL
                            `FUNC_JRL: begin next_state <= `IF; 
                                    r_RegDst<=2; r_MemRead<=0; r_RegWrite<=1;
                                    r_PCSource<=2; r_PCWrite<=1; r_PCWriteCond<=0;
                                    r_Halt<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_OutWrite<=0;
                                    r_next_num_inst <= r_num_inst + 1;
                                    end
                            //WWD
                            `FUNC_WWD: begin next_state <= `IF;
                                    r_OutWrite<=1;
                                    r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_PCWriteCond<=0;
                                    r_next_num_inst <= r_num_inst + 1;
                                    end
                            //HLT, next state = HALT
                            `FUNC_HLT: begin next_state <= `HALT;
                                    r_Halt<=1;
                                    r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0; r_PCWriteCond<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                                    r_next_num_inst <= r_num_inst + 1;
                                    end
                        endcase
                    `OPCODE_ADI: begin next_state <= `ADI_EX; 
                                    r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                    end
                    `OPCODE_ORI: begin next_state <= `ORI_EX; 
                                    r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                    end
                    `OPCODE_LHI: begin next_state <= `LHI_EX; 
                                    r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                    r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                    end
                    //Branch
                    `OPCODE_BNE: begin next_state <= `BNE_EX; 
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                            r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                            end
                    `OPCODE_BEQ: begin next_state <= `BEQ_EX; 
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                            r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                            end
                    `OPCODE_BGZ: begin next_state <= `BGZ_EX; 
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                            r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                            end
                    `OPCODE_BLZ: begin next_state <= `BLZ_EX; 
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                            r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                            end
                    //Jumps
                    `OPCODE_JMP: begin next_state <= `IF; 
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_CAT_TAR;
                            r_PCSource<=0; r_PCWrite<=1; r_PCWriteCond<=0;
                            r_Halt<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                            r_next_num_inst <= r_num_inst + 1;
                            end
                    `OPCODE_JAL: begin next_state <= `IF; 
                            r_RegDst<=2; r_MemtoReg<=0; r_RegWrite<=1;
                            r_ALUSrcA<=0; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_CAT_TAR;
                            r_PCSource<=0; r_PCWrite<=1; r_PCWriteCond<=0;
                            r_Halt<=0; r_MemRead<=0; r_MemWrite<=0;
                            r_IRWrite<=0; r_OutWrite<=0;
                            r_next_num_inst <= r_num_inst + 1;
                            end
                    //JPR, JRL: covered ahead
                    //WWD, HLT: covered ahead
                    //LWD, SWD
                    `OPCODE_LWD: begin next_state <= `LWD_EX; 
                                r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                end
                    `OPCODE_SWD: begin next_state <= `SWD_EX; 
                                r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                                r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                                end
                endcase

            //EX Stage
            //R-type arithmetic
            `ADD_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_ADD;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `SUB_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_SUB;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `AND_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_AND;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `ORR_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_ORR;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `NOT_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_NOT;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `TCP_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_TCP;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `SHL_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_SHL;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `SHR_EX: begin next_state <= `R_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_SHR;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            //I-type arithmetic
            `ADI_EX: begin next_state <= `I_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `ORI_EX: begin next_state <= `I_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ORI;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `LHI_EX: begin next_state <= `I_WB;
                        r_ALUSrcA<=1; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_LHI;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            //Branch
            `BNE_EX: begin next_state <= `IF;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_BNE;
                        r_PCWriteCond<=1; r_PCSource<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            `BEQ_EX: begin next_state <= `IF;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_BEQ;
                        r_PCWriteCond<=1; r_PCSource<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            `BGZ_EX: begin next_state <= `IF;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_BGZ;
                        r_PCWriteCond<=1; r_PCSource<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            `BLZ_EX: begin next_state <= `IF;
                        r_ALUSrcA<=1; r_ALUSrcB<=0; r_ALUOp<=`ALUCODE_BLZ;
                        r_PCWriteCond<=1; r_PCSource<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            //LWD, SWD
            `LWD_EX: begin next_state <= `LWD_MEM;
                        r_ALUSrcA<=1; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            `SWD_EX: begin next_state <= `SWD_MEM;
                        r_ALUSrcA<=1; r_ALUSrcB<=1; r_ALUOp<=`ALUCODE_ADI;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        end
            
            //MEM Stage
            //LWD
            `LWD_MEM: begin next_state <= `LWD_WB;
                        r_IorD<=1; r_MemRead<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemWrite<=0; r_PCWriteCond<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        end
            //SWD
            `SWD_MEM: begin next_state <= `IF;
                        r_IorD<=1; r_MemWrite<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_PCWriteCond<=0;
                        r_IRWrite<=0; r_RegWrite<=0; r_OutWrite<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end

            //WB Stage
            //R-type arithmetic
            `R_WB: begin next_state <= `IF;
                        r_MemtoReg<=0; r_RegDst<=0; r_RegWrite<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            //I-type arithmetic
            `I_WB: begin next_state <= `IF;
                        r_MemtoReg<=0; r_RegDst<=1; r_RegWrite<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
            //LWD
            `LWD_WB: begin next_state <= `IF;
                        r_MemtoReg<=1; r_RegDst<=1; r_RegWrite<=1;
                        r_Halt<=0; r_PCWrite<=0; r_MemRead<=0; r_MemWrite<=0;
                        r_IRWrite<=0; r_OutWrite<=0; r_PCWriteCond<=0;
                        r_next_num_inst <= r_num_inst + 1;
                        end
        endcase
    end

    //Synchronous state transfer (or async. reset)
    always @(posedge clk or negedge reset_n) begin
        //reset logic
        if (~reset_n) begin
            present_state <= `IDLE;
            r_num_inst <= 1;
            r_next_num_inst <= 1;
        end
        else begin
            //State transfer
            present_state <= next_state;
            r_num_inst <= r_next_num_inst;
        end
    end
endmodule